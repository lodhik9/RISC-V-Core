----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Mario Ivanov
-- 
-- Create Date: 08/06/2022 10:37:40 AM
-- Design Name: 
-- Module Name: Adder_TB - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Adder_TB is

end Adder_TB;

architecture Behavioral of Adder_TB is
component Adder is
    Port ( offsetToJump : in STD_LOGIC_VECTOR (31 downto 0);
           programCounter : in STD_LOGIC_VECTOR (31 downto 0);
           resultingProgramCounter : out STD_LOGIC_VECTOR (31 downto 0));
end component;
signal offsetToJump : STD_LOGIC_VECTOR (31 downto 0);
signal programCounter: STD_LOGIC_VECTOR (31 downto 0) := "00100000000000000000000000000000";
signal resultingProgramCounter: STD_LOGIC_VECTOR(31 downto 0);
begin                                                           -- Offset to jump                     Initial program counter            Expected result
offsetToJump <= "00000000000000000000000000000001" after 20 ns, -- 00000000000000000000000000000001 + 00100000000000000000000000000000 = 00100000000000000000000000000001 
                "00000000000000000000000000000011" after 40 ns, -- 00000000000000000000000000000011 + 00100000000000000000000000000001 = 00100000000000000000000000000100
                "00000000000000000000000000000101" after 60 ns, -- 00000000000000000000000000000101 + 00100000000000000000000000000100 = 00100000000000000000000000001001
                "00000000000000000000000000001001" after 80 ns, -- 00000000000000000000000000001001 + 00100000000000000000000000001001 = 00100000000000000000000000010010
                "00000000000000000000000000010001" after 100 ns, -- 00000000000000000000000000010001 + 00100000000000000000000000010010 = 00100000000000000000000000100011
                "00000000000000000000000000100001" after 110 ns, -- 00000000000000000000000000100001 + 00100000000000000000000000100011 = 0100000000000000000000001000100
                "00000000000000000000000001000001" after 130 ns, -- 00000000000000000000000001000001 + 0100000000000000000000001000100 = 0100000000000000000000010000101
                "00000000000000000000000010000001" after 150 ns, -- 00000000000000000000000010000001 + 0100000000000000000000010000101 = 0100000000000000000000100000110
                "00000000000000000000000100000001" after 170 ns, -- 00000000000000000000000100000001 + 0100000000000000000000100000110 = 0100000000000000000001000000111
                "00000000000000000000001000000001" after 190 ns, -- 00000000000000000000001000000001 + 0100000000000000000001000000111 = 0100000000000000000010000001000
                "00000000000000000000010000000001" after 210 ns, -- 00000000000000000000010000000001 + 0100000000000000000010000001000 = 0100000000000000000100000001001
                "00000000000000000000100000000001" after 230 ns, -- 00000000000000000000100000000001 + 0100000000000000000100000001001 = 0100000000000000001000000001010
                "00000000000000000001000000000001" after 250 ns, -- 00000000000000000001000000000001 + 0100000000000000001000000001010 = 0100000000000000010000000001011
                "00000000000000000010000000000001" after 270 ns, -- 00000000000000000010000000000001 + 0100000000000000010000000001011 = 0100000000000000100000000001100
                "00000000000000000100000000000001" after 290 ns, -- 00000000000000000100000000000001 + 0100000000000000100000000001100 = 0100000000000001000000000001101
                "00000000000000001000000000000001" after 310 ns, -- 00000000000000001000000000000001 + 0100000000000001000000000001101 = 0100000000000010000000000001110
                "00000000000000010000000000000001" after 330 ns, -- 00000000000000010000000000000001 + 0100000000000010000000000001110 = 0100000000000100000000000001111
                "00000000000000100000000000000001" after 350 ns, -- 00000000000000100000000000000001 + 0100000000000100000000000001111 = 0100000000001000000000000010000
                "00000000000001000000000000000001" after 370 ns, -- 00000000000001000000000000000001 + 0100000000001000000000000010000 = 0100000000010000000000000010001
                "00000000000010000000000000000001" after 390 ns, -- 00000000000010000000000000000001 + 0100000000010000000000000010001 = 0100000000100000000000000010010
                "00000000000100000000000000000001" after 410 ns, -- 00000000000100000000000000000001 + 0100000000100000000000000010010 = 0100000001000000000000000010011
                "00000000001000000000000000000001" after 430 ns, -- 00000000001000000000000000000001 + 0100000001000000000000000010011 = 0100000010000000000000000010100
                "00000000010000000000000000000001" after 450 ns, -- 00000000010000000000000000000001 + 0100000010000000000000000010100 = 0100000100000000000000000010101
                "00000000100000000000000000000001" after 470 ns, -- 00000000100000000000000000000001 + 0100000100000000000000000010101 = 0100001000000000000000000010110
                "00000001000000000000000000000001" after 490 ns, -- 00000001000000000000000000000001 + 0100001000000000000000000010110 = 0100010000000000000000000010111
                "00000010000000000000000000000001" after 510 ns, -- 00000010000000000000000000000001 + 0100010000000000000000000010111 = 0100100000000000000000000011000
                "00000100000000000000000000000001" after 530 ns, -- 00000100000000000000000000000001 + 0100100000000000000000000011000 = 0101000000000000000000000011001
                "00001000000000000000000000000001" after 550 ns, -- 00001000000000000000000000000001 + 0101000000000000000000000011001 = 0110000000000000000000000011010
                "00010000000000000000000000000001" after 570 ns, -- 00010000000000000000000000000001 + 0110000000000000000000000011010 = 01000000000000000000000000011011
                "00100000000000000000000000000001" after 590 ns, -- 00100000000000000000000000000001 + 01000000000000000000000000011011 = 01100000000000000000000000011100
                "01000000000000000000000000000001" after 610 ns; -- 01000000000000000000000000000001 + 01100000000000000000000000011100 = 010100000000000000000000000011101

        dut : Adder port map(
            offsetToJump => offsetToJump,
            programCounter => programCounter,
            resultingProgramCounter => resultingProgramCounter
        );

end Behavioral;
